`define cos 992981
`define sin 118273

//`define cos 1000000
//`define sin 0

`define bitsize 64
`define bits (`bitsize-1)
`define clk 5
`define chash 2*`clk

